

`timescale 1ns/1ps

import uvm_pkg::*;
`include "uvm_macros.svh"