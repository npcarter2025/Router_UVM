`ifndef PORT_B_SEQUENCER_SVH
`define PORT_B_SEQUENCER_SVH

typedef uvm_sequencer #(port_b_item) port_b_sequencer;

`endif