`ifndef PORT_A_SEQUENCER_SVH
`define PORT_A_SEQUENCER_SVH

typedef uvm_sequencer #(port_a_item) port_a_sequencer;

`endif