`ifndef DISABLE_VSEQ_SVH
`define DISABLE_VSEQ_SVH

class disable_vseq extends uvm_sequence;
    `uvm_object_utils(disable_vseq)


endclass

`endif