`ifndef REG_SEQUENCER_SVH
`define REG_SEQUENCER_SVH

typedef uvm_sequencer #(reg_item) reg_sequencer;

`endif